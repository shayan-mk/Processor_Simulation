library verilog;
use verilog.vl_types.all;
entity CA_Project is
    port(
        pin_name_2      : in     vl_logic;
        pin_name_1      : in     vl_logic;
        pin_name_5      : in     vl_logic
    );
end CA_Project;
