library verilog;
use verilog.vl_types.all;
entity CA_Project_vlg_vec_tst is
end CA_Project_vlg_vec_tst;
